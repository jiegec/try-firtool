module MulAddRecFNToRaw_preMul(
  input  [1:0]  io_op, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  input  [32:0] io_a, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  input  [32:0] io_b, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  input  [32:0] io_c, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [23:0] io_mulAddA, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [23:0] io_mulAddB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [47:0] io_mulAddC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isSigNaNAny, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isNaNAOrB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isInfA, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isZeroA, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isInfB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isZeroB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_signProd, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isNaNC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isInfC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_isZeroC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [9:0]  io_toPostMul_sExpSum, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_doSubMags, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_CIsDominant, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [4:0]  io_toPostMul_CDom_CAlignDist, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output [25:0] io_toPostMul_highAlignedSigC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
  output        io_toPostMul_bit0AlignedSigC // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 73:16]
);
  wire [8:0] rawA_exp = io_a[31:23]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 51:21]
  wire  rawA_isZero = rawA_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  wire  rawA_isSpecial = rawA_exp[8:7] == 2'h3; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 53:53]
  wire  rawA__isNaN = rawA_isSpecial & rawA_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 56:33]
  wire  rawA__sign = io_a[32]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 59:25]
  wire [9:0] rawA__sExp = {1'b0,$signed(rawA_exp)}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 60:27]
  wire  _rawA_out_sig_T = ~rawA_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:35]
  wire [24:0] rawA__sig = {1'h0,_rawA_out_sig_T,io_a[22:0]}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:44]
  wire [8:0] rawB_exp = io_b[31:23]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 51:21]
  wire  rawB_isZero = rawB_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  wire  rawB_isSpecial = rawB_exp[8:7] == 2'h3; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 53:53]
  wire  rawB__isNaN = rawB_isSpecial & rawB_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 56:33]
  wire  rawB__sign = io_b[32]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 59:25]
  wire [9:0] rawB__sExp = {1'b0,$signed(rawB_exp)}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 60:27]
  wire  _rawB_out_sig_T = ~rawB_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:35]
  wire [24:0] rawB__sig = {1'h0,_rawB_out_sig_T,io_b[22:0]}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:44]
  wire [8:0] rawC_exp = io_c[31:23]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 51:21]
  wire  rawC_isZero = rawC_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  wire  rawC_isSpecial = rawC_exp[8:7] == 2'h3; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 53:53]
  wire  rawC__isNaN = rawC_isSpecial & rawC_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 56:33]
  wire  rawC__sign = io_c[32]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 59:25]
  wire [9:0] rawC__sExp = {1'b0,$signed(rawC_exp)}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 60:27]
  wire  _rawC_out_sig_T = ~rawC_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:35]
  wire [24:0] rawC__sig = {1'h0,_rawC_out_sig_T,io_c[22:0]}; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 61:44]
  wire  signProd = rawA__sign ^ rawB__sign ^ io_op[1]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 96:42]
  wire [10:0] _sExpAlignedProd_T = $signed(rawA__sExp) + $signed(rawB__sExp); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 99:19]
  wire [10:0] sExpAlignedProd = $signed(_sExpAlignedProd_T) - 11'she5; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 99:32]
  wire  doSubMags = signProd ^ rawC__sign ^ io_op[0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 101:42]
  wire [10:0] _GEN_0 = {{1{rawC__sExp[9]}},rawC__sExp}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 105:42]
  wire [10:0] sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 105:42]
  wire [9:0] posNatCAlignDist = sNatCAlignDist[9:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 106:42]
  wire  isMinCAlign = rawA_isZero | rawB_isZero | $signed(sNatCAlignDist) < 11'sh0; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 107:50]
  wire  CIsDominant = _rawC_out_sig_T & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 109:23]
  wire [6:0] _CAlignDist_T_2 = posNatCAlignDist < 10'h4a ? posNatCAlignDist[6:0] : 7'h4a; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 113:16]
  wire [6:0] CAlignDist = isMinCAlign ? 7'h0 : _CAlignDist_T_2; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 111:12]
  wire [24:0] _mainAlignedSigC_T = ~rawC__sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 119:25]
  wire [24:0] _mainAlignedSigC_T_1 = doSubMags ? _mainAlignedSigC_T : rawC__sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 119:13]
  wire [52:0] _mainAlignedSigC_T_3 = doSubMags ? 53'h1fffffffffffff : 53'h0; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 119:53]
  wire [77:0] _mainAlignedSigC_T_5 = {_mainAlignedSigC_T_1,_mainAlignedSigC_T_3}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 119:94]
  wire [77:0] mainAlignedSigC = $signed(_mainAlignedSigC_T_5) >>> CAlignDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 119:100]
  wire [26:0] _reduced4CExtra_T = {rawC__sig, 2'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 121:30]
  wire  reduced4CExtra_reducedVec_0 = |_reduced4CExtra_T[3:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_1 = |_reduced4CExtra_T[7:4]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_2 = |_reduced4CExtra_T[11:8]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_3 = |_reduced4CExtra_T[15:12]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_4 = |_reduced4CExtra_T[19:16]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_5 = |_reduced4CExtra_T[23:20]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  reduced4CExtra_reducedVec_6 = |_reduced4CExtra_T[26:24]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 123:57]
  wire [6:0] _reduced4CExtra_T_1 = {reduced4CExtra_reducedVec_6,reduced4CExtra_reducedVec_5,reduced4CExtra_reducedVec_4,
    reduced4CExtra_reducedVec_3,reduced4CExtra_reducedVec_2,reduced4CExtra_reducedVec_1,reduced4CExtra_reducedVec_0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 124:20]
  wire [32:0] reduced4CExtra_shift = 33'sh100000000 >>> CAlignDist[6:2]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 76:56]
  wire [5:0] _reduced4CExtra_T_18 = {reduced4CExtra_shift[14],reduced4CExtra_shift[15],reduced4CExtra_shift[16],
    reduced4CExtra_shift[17],reduced4CExtra_shift[18],reduced4CExtra_shift[19]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [6:0] _GEN_1 = {{1'd0}, _reduced4CExtra_T_18}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 121:68]
  wire [6:0] _reduced4CExtra_T_19 = _reduced4CExtra_T_1 & _GEN_1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 121:68]
  wire  reduced4CExtra = |_reduced4CExtra_T_19; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 129:11]
  wire  _alignedSigC_T_4 = &mainAlignedSigC[2:0] & ~reduced4CExtra; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 133:44]
  wire  _alignedSigC_T_7 = |mainAlignedSigC[2:0] | reduced4CExtra; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 134:44]
  wire  _alignedSigC_T_8 = doSubMags ? _alignedSigC_T_4 : _alignedSigC_T_7; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 132:16]
  wire [74:0] alignedSigC_hi = mainAlignedSigC[77:3]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 131:12]
  wire [75:0] alignedSigC = {alignedSigC_hi,_alignedSigC_T_8}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 131:12]
  wire  _io_toPostMul_isSigNaNAny_T_2 = rawA__isNaN & ~rawA__sig[22]; // @[submodules/berkeley-hardfloat/src/main/scala/common.scala 82:46]
  wire  _io_toPostMul_isSigNaNAny_T_5 = rawB__isNaN & ~rawB__sig[22]; // @[submodules/berkeley-hardfloat/src/main/scala/common.scala 82:46]
  wire  _io_toPostMul_isSigNaNAny_T_9 = rawC__isNaN & ~rawC__sig[22]; // @[submodules/berkeley-hardfloat/src/main/scala/common.scala 82:46]
  wire [10:0] _io_toPostMul_sExpSum_T_2 = $signed(sExpAlignedProd) - 11'sh18; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 157:53]
  wire [10:0] _io_toPostMul_sExpSum_T_3 = CIsDominant ? $signed({{1{rawC__sExp[9]}},rawC__sExp}) : $signed(
    _io_toPostMul_sExpSum_T_2); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 157:12]
  assign io_mulAddA = rawA__sig[23:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 140:16]
  assign io_mulAddB = rawB__sig[23:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 141:16]
  assign io_mulAddC = alignedSigC[48:1]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 142:30]
  assign io_toPostMul_isSigNaNAny = _io_toPostMul_isSigNaNAny_T_2 | _io_toPostMul_isSigNaNAny_T_5 |
    _io_toPostMul_isSigNaNAny_T_9; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 145:58]
  assign io_toPostMul_isNaNAOrB = rawA__isNaN | rawB__isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 147:42]
  assign io_toPostMul_isInfA = rawA_isSpecial & ~rawA_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 57:33]
  assign io_toPostMul_isZeroA = rawA_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  assign io_toPostMul_isInfB = rawB_isSpecial & ~rawB_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 57:33]
  assign io_toPostMul_isZeroB = rawB_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  assign io_toPostMul_signProd = rawA__sign ^ rawB__sign ^ io_op[1]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 96:42]
  assign io_toPostMul_isNaNC = rawC_isSpecial & rawC_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 56:33]
  assign io_toPostMul_isInfC = rawC_isSpecial & ~rawC_exp[6]; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 57:33]
  assign io_toPostMul_isZeroC = rawC_exp[8:6] == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/rawFloatFromRecFN.scala 52:53]
  assign io_toPostMul_sExpSum = _io_toPostMul_sExpSum_T_3[9:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 156:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC__sign ^ io_op[0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 101:42]
  assign io_toPostMul_CIsDominant = _rawC_out_sig_T & (isMinCAlign | posNatCAlignDist <= 10'h18); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 109:23]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[4:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 160:47]
  assign io_toPostMul_highAlignedSigC = alignedSigC[74:49]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 162:20]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 163:48]
endmodule
module MulAddRecFNToRaw_postMul(
  input         io_fromPreMul_isSigNaNAny, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isNaNAOrB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isInfA, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isZeroA, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isInfB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isZeroB, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_signProd, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isNaNC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isInfC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_isZeroC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input  [9:0]  io_fromPreMul_sExpSum, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_doSubMags, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_CIsDominant, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input  [4:0]  io_fromPreMul_CDom_CAlignDist, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input  [25:0] io_fromPreMul_highAlignedSigC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input         io_fromPreMul_bit0AlignedSigC, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input  [48:0] io_mulAddResult, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  input  [2:0]  io_roundingMode, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output        io_invalidExc, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output        io_rawOut_isNaN, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output        io_rawOut_isInf, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output        io_rawOut_isZero, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output        io_rawOut_sign, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output [9:0]  io_rawOut_sExp, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
  output [26:0] io_rawOut_sig // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 170:16]
);
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 184:45]
  wire  opSignC = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 188:42]
  wire [25:0] _sigSum_T_2 = io_fromPreMul_highAlignedSigC + 26'h1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 191:47]
  wire [25:0] _sigSum_T_3 = io_mulAddResult[48] ? _sigSum_T_2 : io_fromPreMul_highAlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 190:16]
  wire [74:0] sigSum = {_sigSum_T_3,io_mulAddResult[47:0],io_fromPreMul_bit0AlignedSigC}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 190:12]
  wire [1:0] _CDom_sExp_T = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 201:69]
  wire [9:0] _GEN_0 = {{8{_CDom_sExp_T[1]}},_CDom_sExp_T}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 201:43]
  wire [9:0] CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 201:43]
  wire [49:0] _CDom_absSigSum_T_1 = ~sigSum[74:25]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 204:13]
  wire [49:0] _CDom_absSigSum_T_5 = {1'h0,io_fromPreMul_highAlignedSigC[25:24],sigSum[72:26]}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 207:71]
  wire [49:0] CDom_absSigSum = io_fromPreMul_doSubMags ? _CDom_absSigSum_T_1 : _CDom_absSigSum_T_5; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 203:12]
  wire [23:0] _CDom_absSigSumExtra_T_1 = ~sigSum[24:1]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 213:14]
  wire  _CDom_absSigSumExtra_T_2 = |_CDom_absSigSumExtra_T_1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 213:36]
  wire  _CDom_absSigSumExtra_T_4 = |sigSum[25:1]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 214:37]
  wire  CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _CDom_absSigSumExtra_T_2 : _CDom_absSigSumExtra_T_4; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 212:12]
  wire [80:0] _GEN_5 = {{31'd0}, CDom_absSigSum}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 217:24]
  wire [80:0] _CDom_mainSig_T = _GEN_5 << io_fromPreMul_CDom_CAlignDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 217:24]
  wire [28:0] CDom_mainSig = _CDom_mainSig_T[49:21]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 217:56]
  wire [26:0] _CDom_reduced4SigExtra_T_1 = {CDom_absSigSum[23:0], 3'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 220:53]
  wire  CDom_reduced4SigExtra_reducedVec_0 = |_CDom_reduced4SigExtra_T_1[3:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_1 = |_CDom_reduced4SigExtra_T_1[7:4]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_2 = |_CDom_reduced4SigExtra_T_1[11:8]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_3 = |_CDom_reduced4SigExtra_T_1[15:12]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_4 = |_CDom_reduced4SigExtra_T_1[19:16]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_5 = |_CDom_reduced4SigExtra_T_1[23:20]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 120:54]
  wire  CDom_reduced4SigExtra_reducedVec_6 = |_CDom_reduced4SigExtra_T_1[26:24]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 123:57]
  wire [6:0] _CDom_reduced4SigExtra_T_2 = {CDom_reduced4SigExtra_reducedVec_6,CDom_reduced4SigExtra_reducedVec_5,
    CDom_reduced4SigExtra_reducedVec_4,CDom_reduced4SigExtra_reducedVec_3,CDom_reduced4SigExtra_reducedVec_2,
    CDom_reduced4SigExtra_reducedVec_1,CDom_reduced4SigExtra_reducedVec_0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 124:20]
  wire [2:0] _CDom_reduced4SigExtra_T_4 = ~io_fromPreMul_CDom_CAlignDist[4:2]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 52:21]
  wire [8:0] CDom_reduced4SigExtra_shift = 9'sh100 >>> _CDom_reduced4SigExtra_T_4; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 76:56]
  wire [5:0] _CDom_reduced4SigExtra_T_20 = {CDom_reduced4SigExtra_shift[1],CDom_reduced4SigExtra_shift[2],
    CDom_reduced4SigExtra_shift[3],CDom_reduced4SigExtra_shift[4],CDom_reduced4SigExtra_shift[5],
    CDom_reduced4SigExtra_shift[6]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [6:0] _GEN_1 = {{1'd0}, _CDom_reduced4SigExtra_T_20}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 220:72]
  wire [6:0] _CDom_reduced4SigExtra_T_21 = _CDom_reduced4SigExtra_T_2 & _GEN_1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 220:72]
  wire  CDom_reduced4SigExtra = |_CDom_reduced4SigExtra_T_21; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 221:73]
  wire  _CDom_sig_T_4 = |CDom_mainSig[2:0] | CDom_reduced4SigExtra | CDom_absSigSumExtra; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 224:61]
  wire [26:0] CDom_sig = {CDom_mainSig[28:3],_CDom_sig_T_4}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 223:12]
  wire  notCDom_signSigSum = sigSum[51]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 230:36]
  wire [50:0] _notCDom_absSigSum_T_1 = ~sigSum[50:0]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 233:13]
  wire [50:0] _GEN_2 = {{50'd0}, io_fromPreMul_doSubMags}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 234:41]
  wire [50:0] _notCDom_absSigSum_T_4 = sigSum[50:0] + _GEN_2; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 234:41]
  wire [50:0] notCDom_absSigSum = notCDom_signSigSum ? _notCDom_absSigSum_T_1 : _notCDom_absSigSum_T_4; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 232:12]
  wire  notCDom_reduced2AbsSigSum_reducedVec_0 = |notCDom_absSigSum[1:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_1 = |notCDom_absSigSum[3:2]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_2 = |notCDom_absSigSum[5:4]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_3 = |notCDom_absSigSum[7:6]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_4 = |notCDom_absSigSum[9:8]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_5 = |notCDom_absSigSum[11:10]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_6 = |notCDom_absSigSum[13:12]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_7 = |notCDom_absSigSum[15:14]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_8 = |notCDom_absSigSum[17:16]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_9 = |notCDom_absSigSum[19:18]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_10 = |notCDom_absSigSum[21:20]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_11 = |notCDom_absSigSum[23:22]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_12 = |notCDom_absSigSum[25:24]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_13 = |notCDom_absSigSum[27:26]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_14 = |notCDom_absSigSum[29:28]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_15 = |notCDom_absSigSum[31:30]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_16 = |notCDom_absSigSum[33:32]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_17 = |notCDom_absSigSum[35:34]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_18 = |notCDom_absSigSum[37:36]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_19 = |notCDom_absSigSum[39:38]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_20 = |notCDom_absSigSum[41:40]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_21 = |notCDom_absSigSum[43:42]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_22 = |notCDom_absSigSum[45:44]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_23 = |notCDom_absSigSum[47:46]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_24 = |notCDom_absSigSum[49:48]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced2AbsSigSum_reducedVec_25 = |notCDom_absSigSum[50]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 106:57]
  wire [5:0] notCDom_reduced2AbsSigSum_lo_lo = {notCDom_reduced2AbsSigSum_reducedVec_5,
    notCDom_reduced2AbsSigSum_reducedVec_4,notCDom_reduced2AbsSigSum_reducedVec_3,notCDom_reduced2AbsSigSum_reducedVec_2
    ,notCDom_reduced2AbsSigSum_reducedVec_1,notCDom_reduced2AbsSigSum_reducedVec_0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 107:20]
  wire [12:0] notCDom_reduced2AbsSigSum_lo = {notCDom_reduced2AbsSigSum_reducedVec_12,
    notCDom_reduced2AbsSigSum_reducedVec_11,notCDom_reduced2AbsSigSum_reducedVec_10,
    notCDom_reduced2AbsSigSum_reducedVec_9,notCDom_reduced2AbsSigSum_reducedVec_8,notCDom_reduced2AbsSigSum_reducedVec_7
    ,notCDom_reduced2AbsSigSum_reducedVec_6,notCDom_reduced2AbsSigSum_lo_lo}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 107:20]
  wire [5:0] notCDom_reduced2AbsSigSum_hi_lo = {notCDom_reduced2AbsSigSum_reducedVec_18,
    notCDom_reduced2AbsSigSum_reducedVec_17,notCDom_reduced2AbsSigSum_reducedVec_16,
    notCDom_reduced2AbsSigSum_reducedVec_15,notCDom_reduced2AbsSigSum_reducedVec_14,
    notCDom_reduced2AbsSigSum_reducedVec_13}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 107:20]
  wire [25:0] notCDom_reduced2AbsSigSum = {notCDom_reduced2AbsSigSum_reducedVec_25,
    notCDom_reduced2AbsSigSum_reducedVec_24,notCDom_reduced2AbsSigSum_reducedVec_23,
    notCDom_reduced2AbsSigSum_reducedVec_22,notCDom_reduced2AbsSigSum_reducedVec_21,
    notCDom_reduced2AbsSigSum_reducedVec_20,notCDom_reduced2AbsSigSum_reducedVec_19,notCDom_reduced2AbsSigSum_hi_lo,
    notCDom_reduced2AbsSigSum_lo}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 107:20]
  wire [4:0] _notCDom_normDistReduced2_T_26 = notCDom_reduced2AbsSigSum[1] ? 5'h18 : 5'h19; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_27 = notCDom_reduced2AbsSigSum[2] ? 5'h17 : _notCDom_normDistReduced2_T_26; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_28 = notCDom_reduced2AbsSigSum[3] ? 5'h16 : _notCDom_normDistReduced2_T_27; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_29 = notCDom_reduced2AbsSigSum[4] ? 5'h15 : _notCDom_normDistReduced2_T_28; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_30 = notCDom_reduced2AbsSigSum[5] ? 5'h14 : _notCDom_normDistReduced2_T_29; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_31 = notCDom_reduced2AbsSigSum[6] ? 5'h13 : _notCDom_normDistReduced2_T_30; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_32 = notCDom_reduced2AbsSigSum[7] ? 5'h12 : _notCDom_normDistReduced2_T_31; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_33 = notCDom_reduced2AbsSigSum[8] ? 5'h11 : _notCDom_normDistReduced2_T_32; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_34 = notCDom_reduced2AbsSigSum[9] ? 5'h10 : _notCDom_normDistReduced2_T_33; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_35 = notCDom_reduced2AbsSigSum[10] ? 5'hf : _notCDom_normDistReduced2_T_34; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_36 = notCDom_reduced2AbsSigSum[11] ? 5'he : _notCDom_normDistReduced2_T_35; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_37 = notCDom_reduced2AbsSigSum[12] ? 5'hd : _notCDom_normDistReduced2_T_36; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_38 = notCDom_reduced2AbsSigSum[13] ? 5'hc : _notCDom_normDistReduced2_T_37; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_39 = notCDom_reduced2AbsSigSum[14] ? 5'hb : _notCDom_normDistReduced2_T_38; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_40 = notCDom_reduced2AbsSigSum[15] ? 5'ha : _notCDom_normDistReduced2_T_39; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_41 = notCDom_reduced2AbsSigSum[16] ? 5'h9 : _notCDom_normDistReduced2_T_40; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_42 = notCDom_reduced2AbsSigSum[17] ? 5'h8 : _notCDom_normDistReduced2_T_41; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_43 = notCDom_reduced2AbsSigSum[18] ? 5'h7 : _notCDom_normDistReduced2_T_42; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_44 = notCDom_reduced2AbsSigSum[19] ? 5'h6 : _notCDom_normDistReduced2_T_43; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_45 = notCDom_reduced2AbsSigSum[20] ? 5'h5 : _notCDom_normDistReduced2_T_44; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_46 = notCDom_reduced2AbsSigSum[21] ? 5'h4 : _notCDom_normDistReduced2_T_45; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_47 = notCDom_reduced2AbsSigSum[22] ? 5'h3 : _notCDom_normDistReduced2_T_46; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_48 = notCDom_reduced2AbsSigSum[23] ? 5'h2 : _notCDom_normDistReduced2_T_47; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] _notCDom_normDistReduced2_T_49 = notCDom_reduced2AbsSigSum[24] ? 5'h1 : _notCDom_normDistReduced2_T_48; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [4:0] notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[25] ? 5'h0 : _notCDom_normDistReduced2_T_49; // @[src/main/scala/chisel3/util/Mux.scala 47:70]
  wire [5:0] notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 238:56]
  wire [6:0] _notCDom_sExp_T = {1'b0,$signed(notCDom_nearNormDist)}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 239:76]
  wire [9:0] _GEN_3 = {{3{_notCDom_sExp_T[6]}},_notCDom_sExp_T}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 239:46]
  wire [9:0] notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_3); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 239:46]
  wire [113:0] _GEN_6 = {{63'd0}, notCDom_absSigSum}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 241:27]
  wire [113:0] _notCDom_mainSig_T = _GEN_6 << notCDom_nearNormDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 241:27]
  wire [28:0] notCDom_mainSig = _notCDom_mainSig_T[51:23]; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 241:50]
  wire  notCDom_reduced4SigExtra_reducedVec_0 = |notCDom_reduced2AbsSigSum[1:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_1 = |notCDom_reduced2AbsSigSum[3:2]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_2 = |notCDom_reduced2AbsSigSum[5:4]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_3 = |notCDom_reduced2AbsSigSum[7:6]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_4 = |notCDom_reduced2AbsSigSum[9:8]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_5 = |notCDom_reduced2AbsSigSum[11:10]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 103:54]
  wire  notCDom_reduced4SigExtra_reducedVec_6 = |notCDom_reduced2AbsSigSum[12]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 106:57]
  wire [6:0] _notCDom_reduced4SigExtra_T_2 = {notCDom_reduced4SigExtra_reducedVec_6,
    notCDom_reduced4SigExtra_reducedVec_5,notCDom_reduced4SigExtra_reducedVec_4,notCDom_reduced4SigExtra_reducedVec_3,
    notCDom_reduced4SigExtra_reducedVec_2,notCDom_reduced4SigExtra_reducedVec_1,notCDom_reduced4SigExtra_reducedVec_0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 107:20]
  wire [3:0] _notCDom_reduced4SigExtra_T_4 = ~notCDom_normDistReduced2[4:1]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 52:21]
  wire [16:0] notCDom_reduced4SigExtra_shift = 17'sh10000 >>> _notCDom_reduced4SigExtra_T_4; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 76:56]
  wire [5:0] _notCDom_reduced4SigExtra_T_20 = {notCDom_reduced4SigExtra_shift[1],notCDom_reduced4SigExtra_shift[2],
    notCDom_reduced4SigExtra_shift[3],notCDom_reduced4SigExtra_shift[4],notCDom_reduced4SigExtra_shift[5],
    notCDom_reduced4SigExtra_shift[6]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [6:0] _GEN_4 = {{1'd0}, _notCDom_reduced4SigExtra_T_20}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 245:78]
  wire [6:0] _notCDom_reduced4SigExtra_T_21 = _notCDom_reduced4SigExtra_T_2 & _GEN_4; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 245:78]
  wire  notCDom_reduced4SigExtra = |_notCDom_reduced4SigExtra_T_21; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 247:11]
  wire  _notCDom_sig_T_3 = |notCDom_mainSig[2:0] | notCDom_reduced4SigExtra; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 250:39]
  wire [26:0] notCDom_sig = {notCDom_mainSig[28:3],_notCDom_sig_T_3}; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 249:12]
  wire  notCDom_completeCancellation = notCDom_sig[26:25] == 2'h0; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 253:50]
  wire  _notCDom_sign_T = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 257:36]
  wire  notCDom_sign = notCDom_completeCancellation ? roundingMode_min : _notCDom_sign_T; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 255:12]
  wire  notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 262:49]
  wire  notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 263:44]
  wire  notNaN_addZeros = (io_fromPreMul_isZeroA | io_fromPreMul_isZeroB) & io_fromPreMul_isZeroC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 265:58]
  wire  _io_invalidExc_T = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 270:31]
  wire  _io_invalidExc_T_1 = io_fromPreMul_isSigNaNAny | _io_invalidExc_T; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 269:35]
  wire  _io_invalidExc_T_2 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 271:32]
  wire  _io_invalidExc_T_3 = _io_invalidExc_T_1 | _io_invalidExc_T_2; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 270:57]
  wire  _io_invalidExc_T_6 = ~io_fromPreMul_isNaNAOrB & notNaN_isInfProd; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 272:36]
  wire  _io_invalidExc_T_7 = _io_invalidExc_T_6 & io_fromPreMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 273:61]
  wire  _io_invalidExc_T_8 = _io_invalidExc_T_7 & io_fromPreMul_doSubMags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 274:35]
  wire  _io_rawOut_isZero_T_1 = ~io_fromPreMul_CIsDominant & notCDom_completeCancellation; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 281:42]
  wire  _io_rawOut_sign_T_1 = io_fromPreMul_isInfC & opSignC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 284:31]
  wire  _io_rawOut_sign_T_2 = notNaN_isInfProd & io_fromPreMul_signProd | _io_rawOut_sign_T_1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 283:54]
  wire  _io_rawOut_sign_T_5 = notNaN_addZeros & ~roundingMode_min & io_fromPreMul_signProd; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 285:48]
  wire  _io_rawOut_sign_T_6 = _io_rawOut_sign_T_5 & opSignC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 286:36]
  wire  _io_rawOut_sign_T_7 = _io_rawOut_sign_T_2 | _io_rawOut_sign_T_6; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 284:43]
  wire  _io_rawOut_sign_T_9 = io_fromPreMul_signProd | opSignC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 288:37]
  wire  _io_rawOut_sign_T_10 = notNaN_addZeros & roundingMode_min & _io_rawOut_sign_T_9; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 287:46]
  wire  _io_rawOut_sign_T_11 = _io_rawOut_sign_T_7 | _io_rawOut_sign_T_10; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 286:48]
  wire  _io_rawOut_sign_T_15 = io_fromPreMul_CIsDominant ? opSignC : notCDom_sign; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 290:17]
  wire  _io_rawOut_sign_T_16 = ~notNaN_isInfOut & ~notNaN_addZeros & _io_rawOut_sign_T_15; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 289:49]
  assign io_invalidExc = _io_invalidExc_T_3 | _io_invalidExc_T_8; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 271:57]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 276:48]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 263:44]
  assign io_rawOut_isZero = notNaN_addZeros | _io_rawOut_isZero_T_1; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 280:25]
  assign io_rawOut_sign = _io_rawOut_sign_T_11 | _io_rawOut_sign_T_16; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 288:50]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 291:26]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 292:25]
endmodule
module RoundAnyRawFNToRecFN(
  input         io_invalidExc, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input         io_in_isNaN, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input         io_in_isInf, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input         io_in_isZero, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input         io_in_sign, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input  [9:0]  io_in_sExp, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input  [26:0] io_in_sig, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input  [2:0]  io_roundingMode, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  input         io_detectTininess, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  output [32:0] io_out, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
  output [4:0]  io_exceptionFlags // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 57:16]
);
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 89:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 91:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 93:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 94:53]
  wire  roundMagUp = roundingMode_min & io_in_sign | roundingMode_max & ~io_in_sign; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 97:42]
  wire  doShiftSigDown1 = io_in_sig[26]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 119:57]
  wire [8:0] _roundMask_T_1 = ~io_in_sExp[8:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 52:21]
  wire  roundMask_msb = _roundMask_T_1[8]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 58:25]
  wire [7:0] roundMask_lsbs = _roundMask_T_1[7:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 59:26]
  wire  roundMask_msb_1 = roundMask_lsbs[7]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 58:25]
  wire [6:0] roundMask_lsbs_1 = roundMask_lsbs[6:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 59:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[6]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 58:25]
  wire [5:0] roundMask_lsbs_2 = roundMask_lsbs_1[5:0]; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 59:26]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> roundMask_lsbs_2; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 76:56]
  wire [15:0] _GEN_0 = {{8'd0}, roundMask_shift[57:50]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_7 = _GEN_0 & 16'hff; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_9 = {roundMask_shift[49:42], 8'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_11 = _roundMask_T_9 & 16'hff00; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _GEN_1 = {{4'd0}, _roundMask_T_12[15:4]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_17 = _GEN_1 & 16'hf0f; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_19 = {_roundMask_T_12[11:0], 4'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_21 = _roundMask_T_19 & 16'hf0f0; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _GEN_2 = {{2'd0}, _roundMask_T_22[15:2]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_27 = _GEN_2 & 16'h3333; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_29 = {_roundMask_T_22[13:0], 2'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_31 = _roundMask_T_29 & 16'hcccc; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _GEN_3 = {{1'd0}, _roundMask_T_32[15:1]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_37 = _GEN_3 & 16'h5555; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_39 = {_roundMask_T_32[14:0], 1'h0}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_41 = _roundMask_T_39 & 16'haaaa; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [15:0] _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [21:0] _roundMask_T_59 = {_roundMask_T_42,roundMask_shift[58],roundMask_shift[59],roundMask_shift[60],
    roundMask_shift[61],roundMask_shift[62],roundMask_shift[63]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [21:0] _roundMask_T_60 = ~_roundMask_T_59; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 73:32]
  wire [21:0] _roundMask_T_61 = roundMask_msb_2 ? 22'h0 : _roundMask_T_60; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 73:21]
  wire [21:0] _roundMask_T_62 = ~_roundMask_T_61; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 73:17]
  wire [24:0] _roundMask_T_63 = {_roundMask_T_62,3'h7}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 68:58]
  wire [2:0] _roundMask_T_70 = {roundMask_shift[0],roundMask_shift[1],roundMask_shift[2]}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 77:20]
  wire [2:0] _roundMask_T_71 = roundMask_msb_2 ? _roundMask_T_70 : 3'h0; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 62:24]
  wire [24:0] _roundMask_T_72 = roundMask_msb_1 ? _roundMask_T_63 : {{22'd0}, _roundMask_T_71}; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 67:24]
  wire [24:0] _roundMask_T_73 = roundMask_msb ? _roundMask_T_72 : 25'h0; // @[submodules/berkeley-hardfloat/src/main/scala/primitives.scala 62:24]
  wire [24:0] _GEN_4 = {{24'd0}, doShiftSigDown1}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 158:23]
  wire [24:0] _roundMask_T_74 = _roundMask_T_73 | _GEN_4; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 158:23]
  wire [26:0] roundMask = {_roundMask_T_74,2'h3}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 158:42]
  wire [27:0] _shiftedRoundMask_T = {1'h0,_roundMask_T_74,2'h3}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 161:41]
  wire [26:0] shiftedRoundMask = _shiftedRoundMask_T[27:1]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 161:53]
  wire [26:0] _roundPosMask_T = ~shiftedRoundMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 162:28]
  wire [26:0] roundPosMask = _roundPosMask_T & roundMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 162:46]
  wire [26:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 163:40]
  wire  roundPosBit = |_roundPosBit_T; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 163:56]
  wire [26:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 164:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 164:62]
  wire  anyRound = roundPosBit | anyRoundExtra; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 165:36]
  wire  _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 168:38]
  wire  _roundIncr_T_1 = (roundingMode_near_even | roundingMode_near_maxMag) & roundPosBit; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 168:67]
  wire  _roundIncr_T_2 = roundMagUp & anyRound; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 170:29]
  wire  roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 169:31]
  wire [26:0] _roundedSig_T = io_in_sig | roundMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 173:32]
  wire [25:0] _roundedSig_T_2 = _roundedSig_T[26:2] + 25'h1; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 173:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 175:30]
  wire [25:0] _roundedSig_T_7 = roundingMode_near_even & roundPosBit & _roundedSig_T_4 ? roundMask[26:1] : 26'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 174:25]
  wire [25:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 174:21]
  wire [25:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 173:57]
  wire [26:0] _roundedSig_T_10 = ~roundMask; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 179:32]
  wire [26:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 179:30]
  wire [25:0] _roundedSig_T_15 = roundingMode_odd & anyRound ? roundPosMask[26:1] : 26'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 180:24]
  wire [25:0] _GEN_5 = {{1'd0}, _roundedSig_T_11[26:2]}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 179:47]
  wire [25:0] _roundedSig_T_16 = _GEN_5 | _roundedSig_T_15; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 179:47]
  wire [25:0] roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 172:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[25:24])}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 184:76]
  wire [9:0] _GEN_6 = {{7{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 184:40]
  wire [10:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_6); // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 184:40]
  wire [8:0] common_expOut = sRoundedExp[8:0]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 186:37]
  wire [22:0] common_fractOut = doShiftSigDown1 ? roundedSig[23:1] : roundedSig[22:0]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 188:16]
  wire [3:0] _common_overflow_T = sRoundedExp[10:7]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 195:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 195:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 11'sh6b; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 199:31]
  wire  unboundedRange_roundPosBit = doShiftSigDown1 ? io_in_sig[2] : io_in_sig[1]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 202:16]
  wire  unboundedRange_anyRound = doShiftSigDown1 & io_in_sig[2] | |io_in_sig[1:0]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 204:49]
  wire  _unboundedRange_roundIncr_T_1 = _roundIncr_T & unboundedRange_roundPosBit; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 206:67]
  wire  _unboundedRange_roundIncr_T_2 = roundMagUp & unboundedRange_anyRound; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 208:29]
  wire  unboundedRange_roundIncr = _unboundedRange_roundIncr_T_1 | _unboundedRange_roundIncr_T_2; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 207:46]
  wire  roundCarry = doShiftSigDown1 ? roundedSig[25] : roundedSig[24]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 210:16]
  wire [1:0] _common_underflow_T = io_in_sExp[9:8]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 219:49]
  wire  _common_underflow_T_5 = doShiftSigDown1 ? roundMask[3] : roundMask[2]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 220:30]
  wire  _common_underflow_T_6 = anyRound & $signed(_common_underflow_T) <= 2'sh0 & _common_underflow_T_5; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 219:72]
  wire  _common_underflow_T_10 = doShiftSigDown1 ? roundMask[4] : roundMask[3]; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 222:39]
  wire  _common_underflow_T_11 = ~_common_underflow_T_10; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 222:34]
  wire  _common_underflow_T_12 = io_detectTininess & _common_underflow_T_11; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 221:77]
  wire  _common_underflow_T_13 = _common_underflow_T_12 & roundCarry; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 225:38]
  wire  _common_underflow_T_15 = _common_underflow_T_13 & roundPosBit & unboundedRange_roundIncr; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 226:60]
  wire  _common_underflow_T_16 = ~_common_underflow_T_15; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 221:27]
  wire  _common_underflow_T_17 = _common_underflow_T_6 & _common_underflow_T_16; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 220:76]
  wire  common_underflow = common_totalUnderflow | _common_underflow_T_17; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 216:40]
  wire  common_inexact = common_totalUnderflow | anyRound; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 229:49]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 234:34]
  wire  commonCase = ~isNaNOut & ~io_in_isInf & ~io_in_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 236:61]
  wire  overflow = commonCase & common_overflow; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 237:32]
  wire  underflow = commonCase & common_underflow; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 238:32]
  wire  inexact = overflow | commonCase & common_inexact; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 239:28]
  wire  overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 242:60]
  wire  pegMinNonzeroMagOut = commonCase & common_totalUnderflow & (roundMagUp | roundingMode_odd); // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 244:45]
  wire  pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 245:39]
  wire  notNaN_isInfOut = io_in_isInf | overflow & overflow_roundMagUp; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 247:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 249:22]
  wire [8:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 9'h1c0 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 252:18]
  wire [8:0] _expOut_T_2 = ~_expOut_T_1; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 252:14]
  wire [8:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 251:24]
  wire [8:0] _expOut_T_5 = pegMinNonzeroMagOut ? 9'h194 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 256:18]
  wire [8:0] _expOut_T_6 = ~_expOut_T_5; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 256:14]
  wire [8:0] _expOut_T_7 = _expOut_T_3 & _expOut_T_6; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 255:17]
  wire [8:0] _expOut_T_8 = pegMaxFiniteMagOut ? 9'h80 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 260:18]
  wire [8:0] _expOut_T_9 = ~_expOut_T_8; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 260:14]
  wire [8:0] _expOut_T_10 = _expOut_T_7 & _expOut_T_9; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 259:17]
  wire [8:0] _expOut_T_11 = notNaN_isInfOut ? 9'h40 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 264:18]
  wire [8:0] _expOut_T_12 = ~_expOut_T_11; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 264:14]
  wire [8:0] _expOut_T_13 = _expOut_T_10 & _expOut_T_12; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 263:17]
  wire [8:0] _expOut_T_14 = pegMinNonzeroMagOut ? 9'h6b : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 268:16]
  wire [8:0] _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 267:18]
  wire [8:0] _expOut_T_16 = pegMaxFiniteMagOut ? 9'h17f : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 272:16]
  wire [8:0] _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 271:15]
  wire [8:0] _expOut_T_18 = notNaN_isInfOut ? 9'h180 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 276:16]
  wire [8:0] _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 275:15]
  wire [8:0] _expOut_T_20 = isNaNOut ? 9'h1c0 : 9'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 277:16]
  wire [8:0] expOut = _expOut_T_19 | _expOut_T_20; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 276:73]
  wire [22:0] _fractOut_T_2 = isNaNOut ? 23'h400000 : 23'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 280:16]
  wire [22:0] _fractOut_T_3 = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 279:12]
  wire [22:0] _fractOut_T_5 = pegMaxFiniteMagOut ? 23'h7fffff : 23'h0; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 283:13]
  wire [22:0] fractOut = _fractOut_T_3 | _fractOut_T_5; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 282:11]
  wire [9:0] _io_out_T = {signOut,expOut}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 285:23]
  wire [3:0] _io_exceptionFlags_T_2 = {io_invalidExc,1'h0,overflow,underflow}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 287:53]
  assign io_out = {_io_out_T,fractOut}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 285:33]
  assign io_exceptionFlags = {_io_exceptionFlags_T_2,inexact}; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 287:66]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input         io_in_isNaN, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input         io_in_isInf, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input         io_in_isZero, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input         io_in_sign, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input  [9:0]  io_in_sExp, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input  [26:0] io_in_sig, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input  [2:0]  io_roundingMode, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  input         io_detectTininess, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  output [32:0] io_out, // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
  output [4:0]  io_exceptionFlags // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 297:16]
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire [9:0] roundAnyRawFNToRecFN_io_in_sExp; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire [26:0] roundAnyRawFNToRecFN_io_in_sig; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire  roundAnyRawFNToRecFN_io_detectTininess; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire [32:0] roundAnyRawFNToRecFN_io_out; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 308:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundAnyRawFNToRecFN_io_detectTininess),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 316:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 317:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 311:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 314:44]
  assign roundAnyRawFNToRecFN_io_detectTininess = io_detectTininess; // @[submodules/berkeley-hardfloat/src/main/scala/RoundAnyRawFNToRecFN.scala 315:44]
endmodule
module MulAddRecFN(
  input  [1:0]  io_op, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  input  [32:0] io_a, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  input  [32:0] io_b, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  input  [32:0] io_c, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  input  [2:0]  io_roundingMode, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  input         io_detectTininess, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  output [32:0] io_out, // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
  output [4:0]  io_exceptionFlags // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 300:16]
);
  wire [1:0] mulAddRecFNToRaw_preMul_io_op; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_a; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_b; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [32:0] mulAddRecFNToRaw_preMul_io_c; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [23:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [47:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [9:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [4:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire [25:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [4:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [25:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [48:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [2:0] mulAddRecFNToRaw_postMul_io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [9:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire [26:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [9:0] roundRawFNToRecFN_io_in_sExp; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [26:0] roundRawFNToRecFN_io_in_sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire  roundRawFNToRecFN_io_detectTininess; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [32:0] roundRawFNToRecFN_io_out; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
  wire [47:0] _mulAddResult_T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 324:45]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 314:15]
    .io_op(mulAddRecFNToRaw_preMul_io_op),
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 316:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_roundingMode(mulAddRecFNToRaw_postMul_io_roundingMode),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 336:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_detectTininess(roundRawFNToRecFN_io_detectTininess),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 342:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 343:23]
  assign mulAddRecFNToRaw_preMul_io_op = io_op; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 318:35]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 319:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 320:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 321:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 328:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _mulAddResult_T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 325:50]
  assign mulAddRecFNToRaw_postMul_io_roundingMode = io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 331:46]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 337:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 339:39]
  assign roundRawFNToRecFN_io_roundingMode = io_roundingMode; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 340:39]
  assign roundRawFNToRecFN_io_detectTininess = io_detectTininess; // @[submodules/berkeley-hardfloat/src/main/scala/MulAddRecFN.scala 341:41]
endmodule
